library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port(clock        : in std_logic;
         address   : in unsigned(6 downto 0);
         data       : out unsigned(15 downto 0)
    );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(15 downto 0);
    constant conteudo_rom : mem := (
        -- caso endereco => conteudo
        0 => "0001011000000101", -- MOV R3, #5
        1 => "0001100000001000", -- MOV R4, #8
        2 => "0001101000000000", -- MOV R5, #0
        3 => "0011101011000000", -- ADD R5, R3
        4 => "0011101100000000", -- ADD R5, R4
        5 => "0001001000000001", -- MOV R1, #1
        6 => "0100101001000000", -- SUB R5, #1
        7 => "0001001000000000", -- MOV R1, #0
        8 => "1111000000010100", -- JMPS 20
        9 => "0000000000000000",
        10 => "0000000000000000",
        11 => "0000000000000000",
        12 => "0000000000000000",
        13 => "0000000000000000",
        14 => "0000000000000000",
        15 => "0000000000000000",
        16 => "0000000000000000",
        17 => "0000000000000000",
        18 => "0000000000000000",
        19 => "0000000000000000",
        20 => "0010011101000000", -- MOV R3, R5
        21 => "1111000000000011", -- JMPS 3
        -- abaixo: casos omissos => (zero em todos os bits)
        others => (others=>'0')
    );
begin
    process(clock)
    begin
        if(rising_edge(clock)) then
            data <= conteudo_rom(to_integer(address));
        end if;
    end process;
end architecture;